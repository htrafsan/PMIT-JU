module hello();
    initial
      $display("hello, I am remon");
endmodule