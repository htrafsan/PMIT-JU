module vlsi(
    input a,
    input b,
    input c, 
    output z
);

assign z = (a)^(b)^(c); 

endmodule